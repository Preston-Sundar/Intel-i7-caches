module Foo(
	input wire x,
	output wire y
);

assign y = x;
endmodule


// wire q, r;
// Foo f(q, r);

// assign q = 0;
// assign q = 1;
// assign q = 0;

// reg o;


// initial begin


// 	// Foo b(q, r);
// 	$display("q = %d", q);
// 	$display("o = %d", o);
// 	$display("r = %d", r);
// 	$finish(1);
// end
